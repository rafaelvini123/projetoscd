library verilog;
use verilog.vl_types.all;
entity BancoRegistrador_vlg_check_tst is
    port(
        rp_data         : in     vl_logic_vector(15 downto 0);
        rq_data         : in     vl_logic_vector(15 downto 0);
        sampler_rx      : in     vl_logic
    );
end BancoRegistrador_vlg_check_tst;
