library verilog;
use verilog.vl_types.all;
entity BancoRegistrador_vlg_vec_tst is
end BancoRegistrador_vlg_vec_tst;
