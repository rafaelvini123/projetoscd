-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Dec 06 11:19:38 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Controlador IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        data : IN STD_LOGIC_VECTOR(15 DOWNTO 0) := "0000000000000000";
        RF_rp_zero : IN STD_LOGIC := '0';
        PC_clr : OUT STD_LOGIC;
        PC_ld : OUT STD_LOGIC;
        IR_ld : OUT STD_LOGIC;
        I_rd : OUT STD_LOGIC;
        D_addr : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        D_rd : OUT STD_LOGIC;
        D_wr : OUT STD_LOGIC;
        RF_s : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        RF_W_addr : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        RF_W_wr : OUT STD_LOGIC;
        RF_Rp_addr : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        RF_Rp_rd : OUT STD_LOGIC;
        RF_Rq_addr : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        RF_Rq_rd : OUT STD_LOGIC;
        alu_s : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        ld_STOI : OUT STD_LOGIC
    );
END Controlador;

ARCHITECTURE BEHAVIOR OF Controlador IS
    TYPE type_fstate IS (Init,Fetch,Decode,Load,Store,Add,Load_constant,Subtract,Jump_if_zero,Jump_zero_jmp,STOI,Store_2,Load_2,Load_3,STOI_2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,data,RF_rp_zero)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Init;
            PC_clr <= '0';
            PC_ld <= '0';
            IR_ld <= '0';
            I_rd <= '0';
            D_addr <= "00000000";
            D_rd <= '0';
            D_wr <= '0';
            RF_s <= "00";
            RF_W_addr <= "0000";
            RF_W_wr <= '0';
            RF_Rp_addr <= "0000";
            RF_Rp_rd <= '0';
            RF_Rq_addr <= "0000";
            RF_Rq_rd <= '0';
            alu_s <= "00";
            ld_STOI <= '0';
        ELSE
            PC_clr <= '0';
            PC_ld <= '0';
            IR_ld <= '0';
            I_rd <= '0';
            D_addr <= "00000000";
            D_rd <= '0';
            D_wr <= '0';
            RF_s <= "00";
            RF_W_addr <= "0000";
            RF_W_wr <= '0';
            RF_Rp_addr <= "0000";
            RF_Rp_rd <= '0';
            RF_Rq_addr <= "0000";
            RF_Rq_rd <= '0';
            alu_s <= "00";
            ld_STOI <= '0';
            CASE fstate IS
                WHEN Init =>
                    reg_fstate <= Fetch;

                    PC_clr <= '1';
                WHEN Fetch =>
                    reg_fstate <= Decode;

                    IR_ld <= '1';

                    I_rd <= '1';
                WHEN Decode =>
                    IF ((data(15 DOWNTO 12) = "0110")) THEN
                        reg_fstate <= STOI;
                    ELSIF ((data(15 DOWNTO 12) = "0001")) THEN
                        reg_fstate <= Store;
                    ELSIF ((data(15 DOWNTO 12) = "0010")) THEN
                        reg_fstate <= Add;
                    ELSIF ((data(15 DOWNTO 12) = "0011")) THEN
                        reg_fstate <= Load_constant;
                    ELSIF ((data(15 DOWNTO 12) = "0100")) THEN
                        reg_fstate <= Subtract;
                    ELSIF ((data(15 DOWNTO 12) = "0101")) THEN
                        reg_fstate <= Jump_if_zero;
                    ELSE
                        reg_fstate <= Load;
                    END IF;
                WHEN Load =>
                    reg_fstate <= Load_2;

                    D_rd <= '1';

                    D_addr <= data(7 DOWNTO 0);
                WHEN Store =>
                    reg_fstate <= Store_2;

                    RF_Rp_addr <= data(11 DOWNTO 8);

                    RF_Rp_rd <= '1';
                WHEN Add =>
                    reg_fstate <= Fetch;

                    alu_s <= "01";

                    RF_W_wr <= '1';

                    RF_Rp_addr <= data(7 DOWNTO 4);

                    RF_W_addr <= data(11 DOWNTO 8);

                    RF_Rq_addr <= data(3 DOWNTO 0);

                    RF_Rq_rd <= '1';

                    RF_s <= "00";

                    RF_Rp_rd <= '1';
                WHEN Load_constant =>
                    reg_fstate <= Fetch;

                    RF_W_wr <= '1';

                    RF_W_addr <= data(11 DOWNTO 8);

                    RF_s <= "10";
                WHEN Subtract =>
                    reg_fstate <= Fetch;

                    alu_s <= "10";

                    RF_W_wr <= '1';

                    RF_Rp_addr <= data(7 DOWNTO 4);

                    RF_W_addr <= data(11 DOWNTO 8);

                    RF_Rq_addr <= data(3 DOWNTO 0);

                    RF_Rq_rd <= '1';

                    RF_s <= "00";

                    RF_Rp_rd <= '1';
                WHEN Jump_if_zero =>
                    IF ((RF_rp_zero = '1')) THEN
                        reg_fstate <= Jump_zero_jmp;
                    ELSIF ((RF_rp_zero = '0')) THEN
                        reg_fstate <= Fetch;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Jump_if_zero;
                    END IF;

                    RF_Rp_addr <= data(11 DOWNTO 8);

                    RF_Rp_rd <= '1';
                WHEN Jump_zero_jmp =>
                    reg_fstate <= Fetch;

                    PC_ld <= '1';
                WHEN STOI =>
                    reg_fstate <= STOI_2;

                    ld_STOI <= '1';

                    RF_Rp_addr <= data(3 DOWNTO 0);

                    RF_Rq_addr <= data(7 DOWNTO 4);

                    RF_Rq_rd <= '1';

                    RF_Rp_rd <= '1';
                WHEN Store_2 =>
                    reg_fstate <= Fetch;

                    D_wr <= '1';

                    D_addr <= data(7 DOWNTO 0);
                WHEN Load_2 =>
                    reg_fstate <= Load_3;

                    RF_s <= "01";
                WHEN Load_3 =>
                    reg_fstate <= Fetch;

                    RF_W_wr <= '1';

                    RF_W_addr <= data(11 DOWNTO 8);
                WHEN STOI_2 =>
                    reg_fstate <= Fetch;

                    ld_STOI <= '1';

                    D_wr <= '1';
                WHEN OTHERS => 
                    PC_clr <= 'X';
                    PC_ld <= 'X';
                    IR_ld <= 'X';
                    I_rd <= 'X';
                    D_addr <= "XXXXXXXX";
                    D_rd <= 'X';
                    D_wr <= 'X';
                    RF_s <= "XX";
                    RF_W_addr <= "XXXX";
                    RF_W_wr <= 'X';
                    RF_Rp_addr <= "XXXX";
                    RF_Rp_rd <= 'X';
                    RF_Rq_addr <= "XXXX";
                    RF_Rq_rd <= 'X';
                    alu_s <= "XX";
                    ld_STOI <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
