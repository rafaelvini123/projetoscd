library verilog;
use verilog.vl_types.all;
entity Memoria_vlg_vec_tst is
end Memoria_vlg_vec_tst;
